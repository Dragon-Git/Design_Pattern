// Bridge pattern in systemverilog